library verilog;
use verilog.vl_types.all;
entity ARM7_TB is
    generic(
        clk_period      : integer := 10
    );
end ARM7_TB;
