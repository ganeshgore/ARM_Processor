`timescale 10ps / 1ps
// SFTUnit(INA(),.INB(),.OPCODE(),.Cin(),.OUT(),.Cout());
module SFTUnit(INA,INB,OPCODE,Cin,OUT,Cout);

input signed [31:0] INA;
input [31:0] INB;
input signed [31:0] OPCODE;
input Cin;
output reg [31:0] OUT;
output reg Cout;

reg [31:0]Data_IN;
wire [31:0]Data_OUT;
reg [4:0]Sel;
wire [3:0]Decode;



barrel32 Shifter(.Data_IN(Data_IN),.Sel(Sel),.Data_OUT(Data_OUT));
I_Decode Shift_I_Decode(.OPCODE(OPCODE),.Dec(Decode));


always@(INA,INB,OPCODE,Cin,Data_OUT,Decode)
	begin
		case(Decode)
		1:OUT = INA;
		2:OUT = INA;
		11:
			begin
				Data_IN = {24'h000000,OPCODE[7:0]};
				Sel = {OPCODE[11:8],1'b0};
				OUT = Data_OUT;	
				Cout = Data_OUT[31];
			end
		7:
			begin
			Data_IN <= {24'h000,INA[7:0]};
			case (OPCODE[6:4])
				3'B000: {Cout,OUT} = INA<<OPCODE[11:7];
				3'B001: {Cout,OUT} = INA<<INB[4:0];
				3'B010: {OUT,Cout} = INA>>OPCODE[11:7];
				3'B011: {OUT,Cout} = INA>>INB[4:0];
				3'B100: {OUT,Cout} = INA>>>OPCODE[11:7];
				3'B101: {OUT,Cout} = INA>>>INB[4:0];
				3'B110: if(OPCODE[11:7] == 5'b00000)
							begin
								Sel = 5'b00001;
								OUT[30:0] = Data_OUT[30:0];
								Cout = Data_OUT[31];
								OUT[31]  = Cin;
							end
						 else
							begin
								Sel = OPCODE[11:7];
								Cout = Data_OUT[31];
								OUT = Data_OUT;
							end
				3'B111: begin 
							Sel = INB[4:0];
							Cout = Data_OUT[31];
							OUT = Data_OUT;
						 end
				3'B001: OUT = INA;
				3'B011: OUT = INA;
				3'B101: OUT = INA;
				3'B111: OUT = INA;
				endcase
			end
		8:begin
			if(OPCODE[25] == 1'b1)
				OUT = INA<<OPCODE[11:4];
			else
				OUT = {OPCODE[11:0],20'b0}>>>20;
			end
		10:OUT <=  OPCODE[23:0]<<2;
		default OUT = 32'bx;
		endcase
		// $display("ShiftUnit:%t\t%h\t%h\t%h\t%h", $time, INA, INB,OPCODE,OUT);
	end

	
endmodule




module barrel32(Data_IN, Sel, Data_OUT);

input   [31:0]    Data_IN;
input   [4:0]     Sel;
output  [31:0]    Data_OUT;

reg     [31:0]    Lvl1 = 0, Lvl2 = 0, Lvl3 = 0; // not really registers, Verilog compliance
wire    [63:0]    Stage1, Stage2;     // wires to simplify FOR loops
integer           i, j;               // loop variables

always @(*) Lvl1 <= Sel[4] ? {Data_IN[15:0], Data_IN[31:16]} : Data_IN; // rotate {0 | 16} bits

assign Stage1 = {Lvl1, Lvl1};    // wraparound a la Verilog

always @(*)    // rotate {0 | 4 | 8 | 12} bits
  case (Sel[3:2])
     2'b00:  Lvl2 <= Stage1[31:0];       // rotate by 0
     2'b01:  for (i=0; i<=31; i=i+1)  Lvl2[i] <= Stage1[i+4];  // rotate by 4
     2'b10:  for (i=0; i<=31; i=i+1)  Lvl2[i] <= Stage1[i+8];  // rotate by 8
     2'b11:  for (i=0; i<=31; i=i+1)  Lvl2[i] <= Stage1[i+12]; // rotate by 12
  endcase

assign Stage2 = {Lvl2, Lvl2};    // wraparound a la Verilog

always @(*)    // rotate {0 | 1 | 2 | 3} bits
  case (Sel[1:0])
     2'b00:  Lvl3 <= Stage2[31:0];       // rotate by 0
     2'b01:  for (j=0; j<=31; j=j+1)  Lvl3[j] <= Stage2[j+1]; // rotate by 1
     2'b10:  for (j=0; j<=31; j=j+1)  Lvl3[j] <= Stage2[j+2]; // rotate by 2
     2'b11:  for (j=0; j<=31; j=j+1)  Lvl3[j] <= Stage2[j+3]; // rotate by 3
  endcase

assign Data_OUT = Lvl3;

endmodule