library verilog;
use verilog.vl_types.all;
entity SFTUnit_TB is
end SFTUnit_TB;
